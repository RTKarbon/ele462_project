* comment for hpsice

vdd 1 0 vdd

.param vdd=1.2V

R1 1 2 1.013843e-07
R2 3 4 1.009806e-07
R3 5 6 1.105636e-07
R4 7 8 1.163129e-07
R5 9 10 1.202099e-07
R6 11 12 1.023943e-07
R7 13 14 1.114067e-07
R8 15 16 1.092288e-07
R9 17 18 1.002147e-07
R10 19 20 1.064602e-07
L1 2 3 1.000000e-09
L2 4 5 1.000000e-09
L3 6 7 1.000000e-09
L4 8 9 1.000000e-09
L5 10 11 1.000000e-09
L6 12 13 1.000000e-09
L7 14 15 1.000000e-09
L8 16 17 1.000000e-09
L9 18 19 1.000000e-09
L10 20 21 1.000000e-09
C1 3 0 9.863462e-08
C2 5 0 9.902890e-08
C3 7 0 9.044564e-08
C4 9 0 8.597499e-08
C5 11 0 8.318781e-08
C6 13 0 9.766169e-08
C7 15 0 8.976117e-08
C8 17 0 9.155097e-08
C9 19 0 9.978576e-08
C10 21 0 9.393179e-08
VSW 1 0 PULSE (0V 1.2V 5us 0.5us 0.5us 4.5us 10us)

* Analysis
.options nomod post
* type
.tran 1ps 50ns

.END
